--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package cnn_types is

    type state is (H_ok, H_nok, V_nok);

end cnn_types;

package body cnn_types is
 
end cnn_types;
