----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity main_cnn is
end main_cnn;

architecture Behavioral of main_cnn is

begin


end Behavioral;

